VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO demux_1_8
  CLASS BLOCK ;
  FOREIGN demux_1_8 ;
  ORIGIN 0.000 0.000 ;
  SIZE 700.000 BY 700.000 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 24.340 10.640 25.940 688.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 177.940 10.640 179.540 688.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 331.540 10.640 333.140 688.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 485.140 10.640 486.740 688.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 638.740 10.640 640.340 688.400 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 30.030 694.380 31.630 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 183.210 694.380 184.810 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 336.390 694.380 337.990 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 489.570 694.380 491.170 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 642.750 694.380 644.350 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 688.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 688.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 688.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 688.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 688.400 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 26.730 694.380 28.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 179.910 694.380 181.510 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 333.090 694.380 334.690 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 486.270 694.380 487.870 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 639.450 694.380 641.050 ;
    END
  END VPWR
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 696.000 367.240 700.000 367.840 ;
    END
  END clk
  PIN i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 418.690 0.000 418.970 4.000 ;
    END
  END i
  PIN o0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 595.790 696.000 596.070 700.000 ;
    END
  END o0
  PIN o1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 442.040 4.000 442.640 ;
    END
  END o1
  PIN o2
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END o2
  PIN o3
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 627.990 0.000 628.270 4.000 ;
    END
  END o3
  PIN o4
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 221.040 4.000 221.640 ;
    END
  END o4
  PIN o5
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 386.490 696.000 386.770 700.000 ;
    END
  END o5
  PIN o6
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 696.000 588.240 700.000 588.840 ;
    END
  END o6
  PIN o7
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 209.390 0.000 209.670 4.000 ;
    END
  END o7
  PIN sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 663.040 4.000 663.640 ;
    END
  END sel[0]
  PIN sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 173.970 696.000 174.250 700.000 ;
    END
  END sel[1]
  PIN sel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 696.000 142.840 700.000 143.440 ;
    END
  END sel[2]
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 694.140 688.245 ;
      LAYER met1 ;
        RECT 0.070 10.640 694.530 688.400 ;
      LAYER met2 ;
        RECT 0.100 695.720 173.690 696.730 ;
        RECT 174.530 695.720 386.210 696.730 ;
        RECT 387.050 695.720 595.510 696.730 ;
        RECT 596.350 695.720 694.510 696.730 ;
        RECT 0.100 4.280 694.510 695.720 ;
        RECT 0.650 4.000 209.110 4.280 ;
        RECT 209.950 4.000 418.410 4.280 ;
        RECT 419.250 4.000 627.710 4.280 ;
        RECT 628.550 4.000 694.510 4.280 ;
      LAYER met3 ;
        RECT 4.000 664.040 696.000 688.325 ;
        RECT 4.400 662.640 696.000 664.040 ;
        RECT 4.000 589.240 696.000 662.640 ;
        RECT 4.000 587.840 695.600 589.240 ;
        RECT 4.000 443.040 696.000 587.840 ;
        RECT 4.400 441.640 696.000 443.040 ;
        RECT 4.000 368.240 696.000 441.640 ;
        RECT 4.000 366.840 695.600 368.240 ;
        RECT 4.000 222.040 696.000 366.840 ;
        RECT 4.400 220.640 696.000 222.040 ;
        RECT 4.000 143.840 696.000 220.640 ;
        RECT 4.000 142.440 695.600 143.840 ;
        RECT 4.000 10.715 696.000 142.440 ;
  END
END demux_1_8
END LIBRARY

